     
d             d       ////  d d           d d        d  d         d   d     



 d    d       d     d     d     d     d       d     d     d   d         d    d      d d           d      d        d             dFFFF d 