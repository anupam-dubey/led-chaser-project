     rd       88,   d      88$    d     888    d    888     d   88 8     d  88 8      d 88         d88  d      d888  d     d888   d    d88$ 8   d   d88, 8    d  d88,       d d88,        dd88,8 d     dd88$8  d    dd88 8  d   dd88 8   d  dd88      d dd88       ddd888 d    ddd888  d   ddd88 8  d  ddd88$ 8   d ddd88,      dddd88,  d   dddd88,8  d  dddd88$8   d dddd88 8   ddddd88 8d  ddddd88   d ddddd88    dddddd888 d dddddd888  ddddddd88$ 8dddddddd88, 8dddddddd88,  dddddddd88,  dddddddd88,8         88,8         88, 8        88, 8dddddddd88,  dddddddd88,  dddddddd88,8         88,8         88, 8        88, 8dddddddd88,  dddddddd88,  dddddddd88,8         88,8         88, 8        88, 8dddddddd88,  dddddddd88,  dddddddd88,8 AAAAAAAA88,8         88, 888, 8        88,  d      d88,   d    d 88,8   d  d  88,8    dd   88, 8   dd   88, 8  d  d  88,   d    d 88,  d      d88,8         88,8         88, 8       88, 8       88,  &       88,  d       88,8 d      88,8 d      88, 8d&      88, 8&d      88,  d     88,  d     88,8  d&     88,8  &d     88, 8 d    88, 8 d    88,    d&    88,    &d    88,8   d    88,8   d   88, 8   d   88, 8   &&   88,     d   88,     d  88,8     d  88,8     d&  88, 8    &d  88, 8    d  88,      d 88,       d 88,8      &d 88,8      d88, 8     d88, 8      d&88        &d88        d888       d888        d88 8       &88 8       88         88          88,8         88,8         88, 8        88, 8