     e
d           d           d           d           d           d           d           d           d           d d         d d        d  d       d   d      d    d     d     d    d      d   d       d  d        d d         ddd        dd d       dd  d      dd   d     dd    d    dd     d   dd      d  dd       d dd        dddd       ddd d      ddd  d     ddd   d    ddd    d   ddd     d  ddd      d ddd       ddddd      dddd d     dddd  d    dddd   d   dddd    d  dddd     d dddd      dddddd     ddddd d    ddddd  d   ddddd   d  ddddd    d ddddd     ddddddd    dddddd d   dddddd  d  dddddd   d dddddd    dddddddd   ddddddd d  ddddddd  d ddddddd   ddddddddd  dddddddd d dddddddd  dddddddddd ddddddddd ddddddddddddddddddddddddddddddddddddddddddd                                 ddddddddddddddddddddddddddddddddd                                 ddddddddddddddddddddddddddddddddd                                 ddddddddddddddddddddddddddddddddd:::::::::::           d         d d       d   d     d     d   d       d d         d         d d       d   d     d     d   d       d d         d