     T d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d                                d1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@Kd                         1@K                          1@                           1                                                                                                                      d      d      d      d      d    d    d d    d d    d d    d d    d  d   d  d   d  d   d  d   d    dd     dd     dd     dd     d   dd     dd     dd     dd     d  d  d   d  d   d  d   d  d   d  d    d d    d d    d d    d d        d      d      d         d      d      d         d      d      d                           ////////                        >>>>>>>>      d      d      d   RRRRRRRR      d      d      d   >>>>>>>>                        ////////                              d      d      d         d      d      d                                                   