     *
d  d              d   d              d   d             d    d             d    d            d     d         d        d        d         d        d         d       d          d       d          d      d           d   d              d  d               d  d               d d d             d  d d           d   d  d         d  d     d       d   d      d     d     d      d   d      d       d d        d       d         d      d d      d       d   d     d      d     d     d    d       d    d   d         d    d d           d   dd             dd                 d                  d                 d ddddddddddddddd  dddddddddddddddd  ddddddddddddddddd  dddddddddddddddd  444444444444444 d  d   d                 d               