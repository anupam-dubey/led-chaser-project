     �
d        d        d        d        d        d        d        dd      d d     d  d    d   d   d    d  d     d d      dd      ddd     dd d    dd  d   dd   d  dd    d dd     dddd    ddd d   ddd  d  ddd   d ddd    ddddd   dddd d  dddd  d dddd   dddddd  ddddd d ddddd  ddddddd dddddd ddddddddddddddddddddddddddddddddddddddddddddddd                        dddddddddddddddddddddddd                        dddddddddddddddddddddddd                        dddddddddddddddddddddddd66666666        d      d d    d   d  d     dd      dd     d  d   d    d d      d                              %       %       d       d       d      %%      %      d       d       d       d      d      %%      %      d       d       d      d      %%      %      d       d       d       d      d      %%      %      d       d       d       d      d      %%      %      d       d       d       d      d      %%      %      d       d       d       d      d      %%      %      d       d       d       d       d       %                      