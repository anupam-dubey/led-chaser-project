     
P"""""""""ddd"P""""""""ddd""P"""""""ddd"""P""""""ddd""""P"""""ddd"""""P""""ddd""""""P"""ddd"""""""P""ddd""""""""P"ddd"""""""""Pddd