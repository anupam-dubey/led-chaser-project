       d d d d d d d d d d              d d d d d d d d d                d d d d d d d d                  d d d d d d d                    d d d d d d                      d d d d d                        d d d d                          d d d                            d d                              d                              d d                            d d d                          d d d d                        d d d d d                      d d d d d d                    d d d d d d d                  d d d d d d d d                d d d d d d d d d              d d d d d d d d d d            